# v-codes
To design NOT gate circuit
module notgate(a,z);
input a;
output z;
assign z=!a;
endmodule
