/*To design XNOR gate circuit*/
module xnorgate(a,b,z);
  input a,b;
  output z;
  assign z=~(a^b);
endmodule
