/*To design OR gate circuit*/
module orgate(a,b,z);
  input a,b;
  output z;
  assign z=a|b;
endmodule
