/*To design XOR gate circuit*/
module xorgate(a,b,z);
  input a,b;
  output z;
  assign z=a^b;
endmodule
